
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_unsigned.ALL;
use IEEE.STD_LOGIC_arith.ALL;


entity gaussina_fn is
    Port ( A : in STD_LOGIC_VECTOR (15 downto 0);   --input Q6.10 signed
           en : in STD_LOGIC;
           Y : out STD_LOGIC_VECTOR (15 downto 0)); --output Q6.10 signed
end gaussina_fn;

architecture Behavioral of gaussina_fn is

signal D :  STD_LOGIC_VECTOR (15 downto 0):=(others=>'0');
signal D_tem :  STD_LOGIC_VECTOR (15 downto 0):=(others=>'0');

constant sigrsq:integer:=50;
begin
D<= A when A(15)='0' else not(A)+1;
D_tem<="0000000100000000" when D <= "0000000000000000" else
"0000000011111111" when D <= "0000000000000101" else
"0000000011111111" when D <= "0000000000001010" else
"0000000011111111" when D <= "0000000000001111" else
"0000000011111111" when D <= "0000000000010100" else
"0000000011111110" when D <= "0000000000011001" else
"0000000011111110" when D <= "0000000000011110" else
"0000000011111101" when D <= "0000000000100011" else
"0000000011111100" when D <= "0000000000101000" else
"0000000011111011" when D <= "0000000000101110" else
"0000000011111010" when D <= "0000000000110011" else
"0000000011111001" when D <= "0000000000111000" else
"0000000011111000" when D <= "0000000000111101" else
"0000000011110111" when D <= "0000000001000010" else
"0000000011110110" when D <= "0000000001000111" else
"0000000011110100" when D <= "0000000001001100" else
"0000000011110011" when D <= "0000000001010001" else
"0000000011110001" when D <= "0000000001010111" else
"0000000011101111" when D <= "0000000001011100" else
"0000000011101110" when D <= "0000000001100001" else
"0000000011101100" when D <= "0000000001100110" else
"0000000011101010" when D <= "0000000001101011" else
"0000000011101000" when D <= "0000000001110000" else
"0000000011100110" when D <= "0000000001110101" else
"0000000011100100" when D <= "0000000001111010" else
"0000000011100001" when D <= "0000000010000000" else
"0000000011011111" when D <= "0000000010000101" else
"0000000011011101" when D <= "0000000010001010" else
"0000000011011010" when D <= "0000000010001111" else
"0000000011011000" when D <= "0000000010010100" else
"0000000011010101" when D <= "0000000010011001" else
"0000000011010011" when D <= "0000000010011110" else
"0000000011010000" when D <= "0000000010100011" else
"0000000011001101" when D <= "0000000010101000" else
"0000000011001011" when D <= "0000000010101110" else
"0000000011001000" when D <= "0000000010110011" else
"0000000011000101" when D <= "0000000010111000" else
"0000000011000010" when D <= "0000000010111101" else
"0000000010111111" when D <= "0000000011000010" else
"0000000010111100" when D <= "0000000011000111" else
"0000000010111001" when D <= "0000000011001100" else
"0000000010110110" when D <= "0000000011010001" else
"0000000010110011" when D <= "0000000011010111" else
"0000000010110000" when D <= "0000000011011100" else
"0000000010101101" when D <= "0000000011100001" else
"0000000010101010" when D <= "0000000011100110" else
"0000000010100111" when D <= "0000000011101011" else
"0000000010100100" when D <= "0000000011110000" else
"0000000010100001" when D <= "0000000011110101" else
"0000000010011110" when D <= "0000000011111010" else
"0000000010011011" when D <= "0000000100000000" else
"0000000010011000" when D <= "0000000100000101" else
"0000000010010101" when D <= "0000000100001010" else
"0000000010010001" when D <= "0000000100001111" else
"0000000010001110" when D <= "0000000100010100" else
"0000000010001011" when D <= "0000000100011001" else
"0000000010001000" when D <= "0000000100011110" else
"0000000010000101" when D <= "0000000100100011" else
"0000000010000010" when D <= "0000000100101000" else
"0000000001111111" when D <= "0000000100101110" else
"0000000001111100" when D <= "0000000100110011" else
"0000000001111001" when D <= "0000000100111000" else
"0000000001110110" when D <= "0000000100111101" else
"0000000001110011" when D <= "0000000101000010" else
"0000000001110000" when D <= "0000000101000111" else
"0000000001101101" when D <= "0000000101001100" else
"0000000001101011" when D <= "0000000101010001" else
"0000000001101000" when D <= "0000000101010111" else
"0000000001100101" when D <= "0000000101011100" else
"0000000001100010" when D <= "0000000101100001" else
"0000000001100000" when D <= "0000000101100110" else
"0000000001011101" when D <= "0000000101101011" else
"0000000001011010" when D <= "0000000101110000" else
"0000000001011000" when D <= "0000000101110101" else
"0000000001010101" when D <= "0000000101111010" else
"0000000001010011" when D <= "0000000110000000" else
"0000000001010000" when D <= "0000000110000101" else
"0000000001001110" when D <= "0000000110001010" else
"0000000001001011" when D <= "0000000110001111" else
"0000000001001001" when D <= "0000000110010100" else
"0000000001000111" when D <= "0000000110011001" else
"0000000001000100" when D <= "0000000110011110" else
"0000000001000010" when D <= "0000000110100011" else
"0000000001000000" when D <= "0000000110101000" else
"0000000000111110" when D <= "0000000110101110" else
"0000000000111100" when D <= "0000000110110011" else
"0000000000111010" when D <= "0000000110111000" else
"0000000000111000" when D <= "0000000110111101" else
"0000000000110110" when D <= "0000000111000010" else
"0000000000110100" when D <= "0000000111000111" else
"0000000000110010" when D <= "0000000111001100" else
"0000000000110000" when D <= "0000000111010001" else
"0000000000101111" when D <= "0000000111010111" else
"0000000000101101" when D <= "0000000111011100" else
"0000000000101011" when D <= "0000000111100001" else
"0000000000101010" when D <= "0000000111100110" else
"0000000000101000" when D <= "0000000111101011" else
"0000000000100110" when D <= "0000000111110000" else
"0000000000100101" when D <= "0000000111110101" else
"0000000000100100" when D <= "0000000111111010" else
"0000000000100010" when D <= "0000001000000000" else
"0000000000100001" when D <= "0000001000000101" else
"0000000000011111" when D <= "0000001000001010" else
"0000000000011110" when D <= "0000001000001111" else
"0000000000011101" when D <= "0000001000010100" else
"0000000000011100" when D <= "0000001000011001" else
"0000000000011011" when D <= "0000001000011110" else
"0000000000011001" when D <= "0000001000100011" else
"0000000000011000" when D <= "0000001000101000" else
"0000000000010111" when D <= "0000001000101110" else
"0000000000010110" when D <= "0000001000110011" else
"0000000000010101" when D <= "0000001000111000" else
"0000000000010100" when D <= "0000001000111101" else
"0000000000010011" when D <= "0000001001000010" else
"0000000000010011" when D <= "0000001001000111" else
"0000000000010010" when D <= "0000001001001100" else
"0000000000010001" when D <= "0000001001010001" else
"0000000000010000" when D <= "0000001001010111" else
"0000000000001111" when D <= "0000001001011100" else
"0000000000001111" when D <= "0000001001100001" else
"0000000000001110" when D <= "0000001001100110" else
"0000000000001101" when D <= "0000001001101011" else
"0000000000001101" when D <= "0000001001110000" else
"0000000000001100" when D <= "0000001001110101" else
"0000000000001011" when D <= "0000001001111010" else
"0000000000001011" when D <= "0000001010000000" else
"0000000000001010" when D <= "0000001010000101" else
"0000000000001010" when D <= "0000001010001010" else
"0000000000000000" ;
Y<=D_tem when en='1';
end Behavioral;
